    // DDR4
    output [0:0]  c0_ddr4_act_n         ,
    output [16:0] c0_ddr4_adr           ,
    output [1:0]  c0_ddr4_ba            ,
    output [1:0]  c0_ddr4_bg            ,
    output [0:0]  c0_ddr4_ck_c          ,
    output [0:0]  c0_ddr4_ck_t          ,
    output [0:0]  c0_ddr4_cke           ,
    output [0:0]  c0_ddr4_cs_n          ,
    inout  [71:0] c0_ddr4_dq            ,
    inout  [17:0] c0_ddr4_dqs_c         ,
    inout  [17:0] c0_ddr4_dqs_t         ,
    output [0:0]  c0_ddr4_odt           ,
    output [0:0]  c0_ddr4_par           ,
    output [0:0]  c0_ddr4_reset_n       ,
