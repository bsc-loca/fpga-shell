    // CMS
    input [0:0]   satellite_uart_rxd    ,
    output [0:0]  satellite_uart_txd    ,
    input [3:0]   satellite_gpio        ,
    